module hazard_unit(
    input [1:0] reg_wr_ctrl_IDEX,       //Is instruction in EX stage a load instruction?
    input [`REG_FIELD_RANGE] rd_IDEX,   //what register will EX stage instruction load to?

    input [`REG_FIELD_RANGE] rs1_ID, rs2_ID,    //what source registers are we using in ID?
    input pc_rs1_sel, imm_rs2_sel,             //Are these fields of the ID instruction truly register addresses?
);

endmodule