module MMM_wrapper #(
    parameter  INW              = 32,
    parameter  OUTW             = 32,
    parameter  M                = 16,
    parameter  N                = 16,
    parameter  MAXK             = 16,
    localparam K_BITS           = $clog2(MAXK+1),
    localparam A_ADDR_BITS      = $clog2(M*MAXK),
    localparam B_ADDR_BITS      = $clog2(MAXK*N),
    localparam OUT_ADDR_BITS    = $clog2(M*N)
)(
    input clk, reset,

    input [INW-1:0] K_in,   //remember to add a flipflop for K value
    input start_mmm,        //generated by that set/clr flipflop
    input wait_mmm_finish,

    input [INW-1:0]  mata_data, matb_data,
    output logic [A_ADDR_BITS-1:0] mata_rdaddr,
    output logic [B_ADDR_BITS-1:0] matb_rdaddr,

    output logic [INW-1:0] outmat_data,             
    output logic [OUT_ADDR_BITS-1:0] outmat_wraddr,  //delay the address, and wren by 1 cycle because of pipeline
    output logic outmat_wren,

    output logic stall       
);

    logic compute_start, compute_finished;
    logic [K_BITS-1:0] new_K;
    always_ff @(posedge clk) begin
        if(reset) begin
            compute_start <= 0;
        end
        else begin
            if(start_mmm) 
                compute_start <= 1;
            else if(compute_finished)
                compute_start <= 0;
        end
    end

    always_ff @(posedge clk) begin
        if(reset)
            new_K <= 0;
        else
            new_K <= K_in[K_BITS-1:0];
    end

    MMM #(.INW(INW), .OUTW(OUTW), .M(M), .N(N), .MAXK(MAXK)) MMM (.*);

    assign stall = (compute_start & wait_mmm_finish);

endmodule