`include "inst_defs.sv"
